--Processador
--PC
--Bibliotecas e pacotes
LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
--Entidade
entity Processador is
	port(
	
	);
end entity;	
architecture Behavior of Processador is
begin
	
end architecture;