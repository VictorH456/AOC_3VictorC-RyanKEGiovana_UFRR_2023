--Ram
--Bibliotecas e pacotes
LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
--Entidade
entity Ram is
	port(
	
	);
end entity;	
architecture Behavior of Ram is
begin
	
end architecture;