--Ula
--Bibliotecas e pacotes
LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
--Entidade
entity Ula is

end entity;
architecture Behavior of ula is
begin
	
end architecture;