--Unidade de controle
--Bibliotecas e pacotes
LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
--Entidade
entity Uc is

end entity;
architecture Behavior of Uc is
begin
	
end architecture;