--Registradores
--Bibliotecas e pacotes
LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
--Entidade
entity PC is
	port(
	
	);
end entity;	
architecture Behavior of Registradores is
begin
	
end architecture;