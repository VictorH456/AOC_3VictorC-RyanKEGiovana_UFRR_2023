  LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

Entity REGISTRADORES is 
	port(
	Clock, Reg_Write: IN STD_LOGIC;
	Reg1: IN STD_LOGIC_VECTOR (3 DOWNTO 0); -- nomeclatura do vetor
	Reg2: IN STD_LOGIC_VECTOR (3 DOWNTO 0); -- nomeclatura do vetor
	Reg3: IN STD_LOGIC_VECTOR (3 DOWNTO 0); -- nomeclatura do vetor
	Write_data: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
	RegA_de_saida: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
	RegB_de_saida: OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
	);
END REGISTRADORES;
ARCHITECTURE BEHAVIOR OF REGISTRADORES IS
TYPE REGISTRADORES IS ARRAY (0 TO 8) OF STD_LOGIC_VECTOR (15 DOWNTO 0);
SIGNAL MEM_REGISTRADORES: REGISTRADORES;
BEGIN
	PROCESS(Clock, Reg1, Reg2)
	BEGIN
		IF RISING_EDGE(Clock) THEN
			IF (Reg_Write = '1') THEN
				MEM_REGISTRADORES(TO_INTEGER(UNSIGNED(Reg1))) <= Write_data;
			END IF;
		END IF;
		RegA_de_saida <= MEM_REGISTRADORES(TO_INTEGER(UNSIGNED(Reg2))); 
		RegB_de_saida <= MEM_REGISTRADORES(TO_INTEGER(UNSIGNED(Reg3)));
	END PROCESS;
END architecture;	