--Rom
--Bibliotecas e pacotes
LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
--Entidade
entity Rom is
	port(
	
	);
end entity;	
architecture Behavior of Rom is
begin
	
end architecture;